`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// _CPUSystemany: 
// Engineer: 
// 
// Create Date: 21.05.2022 12:52:19
// Design Name: 
// Module Name: sim
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module Project1Test();
    //Input Registers of ALUSystem
    reg[2:0] RF_O1Sel; 
    reg[2:0] RF_O2Sel; 
    reg[1:0] RF_FunSel;
    reg[3:0] RF_RSel;
    reg[3:0] RF_TSel;
    reg[3:0] ALU_FunSel;
    reg[1:0] ARF_OutASel; 
    reg[1:0] ARF_OutBSel; 
    reg[1:0] ARF_FunSel;
    reg[3:0] ARF_RSel;
    reg      IR_LH;
    reg      IR_Enable;
    reg[1:0]      IR_Funsel;
    reg      Mem_WR;
    reg      Mem_CS;
    reg[1:0] MuxASel;
    reg[1:0] MuxBSel;
    reg MuxCSel;
    reg      Clock;
    
    //Test Bench Connection of ALU System
    ALUSystem _ALUSystem(
        .RF_O1Sel(RF_O1Sel), 
        .RF_O2Sel(RF_O2Sel), 
        .RF_FunSel(RF_FunSel),
        .RF_RSel(RF_RSel),
        .RF_TSel(RF_TSel),
        .ALU_FunSel(ALU_FunSel),
        .ARF_OutASel(ARF_OutASel), 
        .ARF_OutBSel(ARF_OutBSel), 
        .ARF_FunSel(ARF_FunSel),
        .ARF_RegSel(ARF_RSel),
        .IR_LH(IR_LH),
        .IR_Enable(IR_Enable),
        .IR_Funsel(IR_Funsel),
        .Mem_WR(Mem_WR),
        .Mem_CS(Mem_CS),
        .MuxASel(MuxASel),
        .MuxBSel(MuxBSel),
        .MuxCSel(MuxCSel),
        .Clock(Clock)
        );
    
    //Test Vector Variables
    reg [41:0] VectorNum, Errors, TotalLine; 
    reg [41:0] TestVectors[3:0];
    reg Reset, Operation;
    initial begin
        Reset = 0;
    end
    //Clock Signal Generation
    always 
    begin
        Clock = 1; #5; Clock = 0; #5; // 10ns period
    end
    
    //Read Test Bench Values
    initial begin
        $readmemb("TestBench.mem", TestVectors); // Read vectors
        VectorNum = 0; Errors = 0; TotalLine=0; Reset=0;// Initialize
    end
    
    // Apply test vectors on rising edge of clock
    always @(posedge Clock)
    begin
        #1; 
        {Operation, RF_O1Sel, RF_O2Sel, RF_FunSel, 
        RF_RSel, RF_TSel, ALU_FunSel, ARF_OutASel, ARF_OutBSel, 
        ARF_FunSel, ARF_RSel, IR_LH, IR_Enable, IR_Funsel, 
        Mem_WR, Mem_CS, MuxASel, MuxBSel, MuxCSel} = TestVectors[VectorNum];
    end
    
    // Check results on falling edge of clk
    always @(negedge Clock)
        if (~Reset) // skip during reset
        begin
            $display("Input Values:");
            $display("Operation: %d", Operation);
            $display("Register File: O1Sel: %d, O2Sel: %d, FunSel: %d, RSel: %d, TSel: %d", RF_O1Sel, RF_O2Sel, RF_FunSel, RF_RSel, RF_TSel);            
            $display("ALU FunSel: %d", ALU_FunSel);
            $display("Addres Register File: OutASel: %d, OutBSel: %d, FunSel: %d, Regsel: %d", ARF_OutASel, ARF_OutBSel, ARF_FunSel, ARF_RSel);            
            $display("Instruction Register: LH: %d, Enable: %d, FunSel: %d", IR_LH, IR_Enable, IR_Funsel);            
            $display("Memory: WR: %d, CS: %d", Mem_WR, Mem_CS);
            $display("MuxASel: %d, MuxBSel: %d, MuxCSel: %d", MuxASel, MuxBSel, MuxCSel);
            
            $display("");
            $display("Output Values:");
            $display("Register File: AOut: %d, BOut: %d", _ALUSystem.AOut, _ALUSystem.BOut);            
            $display("ALUOut: %d, ALUOutFlag: %d, ALUOutFlags: Z:%d, C:%d, N:%d, O:%d,", _ALUSystem.ALUOut, _ALUSystem.ALUOutFlag, _ALUSystem.ALUOutFlag[3],_ALUSystem.ALUOutFlag[2],_ALUSystem.ALUOutFlag[1],_ALUSystem.ALUOutFlag[0]);
            $display("Address Register File: AOut: %d, BOut (Address): %d", _ALUSystem.AOut, _ALUSystem.Address);            
            $display("Memory Out: %d", _ALUSystem.MemoryOut);            
            $display("Instruction Register: IROut: %d", _ALUSystem.IROut);            
            $display("MuxAOut: %d, MuxBOut: %d, MuxCOut: %d", _ALUSystem.MuxAOut, _ALUSystem.MuxBOut, _ALUSystem.MuxCOut);
            
            // increment array index and read next testvector
            VectorNum = VectorNum + 1;
            if (TestVectors[VectorNum] === 42'bx)
            begin
                $display("%d tests completed.",
                VectorNum);
                $finish; // End simulation
            end
        end
endmodule


module Project2Test();
    reg Clock, Reset;
    reg [7:0] T;
    
    always 
        begin
            Clock = 1; #5; Clock = 0; #5; // 10ns period
        end
        
        //reset at start
        initial 
        begin
            Reset = 1; #10; Reset = 0;
        end
        
        initial begin
           // T = 8'h0; #10; T = 8'h1;#10;T = 8'h2;#10T = 8'h3;#10;T = 8'h4;#10;
           T = 8'h0; #10;
        end
    
    always 
    begin
        Clock = 1; #5; Clock = 0; #5; // 10ns period
    end
    
    initial
    begin
       #250; $finish; //this may change
    end
    
    always @(posedge Clock)
        begin
            #10;
            $display("");
            $display("");
            
            $display("input");
            $display("Register File: OutASel: %d, OutBSel: %d, FunSel: %b, Regsel: %b", _CPUSystem.RF_O1Sel, _CPUSystem.RF_O2Sel, _CPUSystem.RF_FunSel, _CPUSystem.RF_RSel);            
            $display("ALU FunSel: %b", _CPUSystem.ALU_FunSel);
            $display("Addres Register File: OutCSel: %d, OutDSel: %d, FunSel: %b, Regsel: %b", _CPUSystem.ARF_OutASel, _CPUSystem.ARF_OutBSel, _CPUSystem.ARF_FunSel, _CPUSystem.ARF_RegSel);            
            $display("Instruction Register: LH: %d, Enable: %d, FunSel: %b", _CPUSystem.IR_LH, _CPUSystem.IR_Enable, _CPUSystem.IR_Funsel);            
            $display("Memory: WR: %d, CS: %d", _CPUSystem.Mem_WR, _CPUSystem.Mem_CS);
            $display("MuxASel: %b, MuxBSel: %b, MuxCSel: %b", _CPUSystem.MuxASel, _CPUSystem.MuxBSel, _CPUSystem.MuxCSel);
            
            $display("");
            $display("output");
            $display("Register File: AOut: %d, BOut: %d", _CPUSystem.ALU_System.AOut, _CPUSystem.ALU_System.BOut);            
            $display("ALUOut: %d, ALUOutFlag: %b, ALUOutFlags: Z:%d, C:%d, N:%d, O:%d,", _CPUSystem.ALU_System.ALUOut, _CPUSystem.ALU_System.ALUOutFlag, _CPUSystem.ALU_System.ALUOutFlag[3],_CPUSystem.ALU_System.ALUOutFlag[2],_CPUSystem.ALU_System.ALUOutFlag[1],_CPUSystem.ALU_System.ALUOutFlag[0]);
            $display("Address Register File: COut: %d, DOut (Address): %d", _CPUSystem.ALU_System.ARF_AOut, _CPUSystem.ALU_System.Address);            
            $display("Memory Out: %d", _CPUSystem.ALU_System.MemoryOut);            
            $display("IROut: %h", _CPUSystem.ALU_System.IROut);
            $display("MuxAOut: %d, MuxBOut: %d, MuxCOut: %d", _CPUSystem.ALU_System.MuxAOut, _CPUSystem.ALU_System.MuxBOut, _CPUSystem.ALU_System.MuxCOut);
                    
        end
    
    CPUSystem _CPUSystem( 
            .Clock(Clock),
            .Reset(Reset),
            .T(T)    
        );
endmodule

